library IEEE;
use IEEE.std_logic_1164.all;
use WORK.myTypes.all;

entity tb_ALU is 
end entity;

architecture test of tb_ALU is 

	component ALU
	generic(NBIT: integer:=32);
	port(
	 	A,B: in std_logic_vector(NBIT-1 downto 0);		
		FUNC: in aluOp;											
		ALU_OUT: out std_logic_vector(31 downto 0);
		OVF: out std_logic);
	end component;
	
	constant clk_period: time := 1 ns;
	signal in_A: std_logic_vector(31 downto 0);
	signal in_B: std_logic_vector(31 downto 0);
	signal op: aluOp;
	signal output: std_logic_vector(31 downto 0);
	signal ovf: std_logic;
	
	begin
	
	ALU1: ALU port map (in_A, in_B, op, output, ovf);
	
		test_proc: process
			begin
			
			in_A <= "00000000000000000000000000001010"; -- 10
			in_B <= "00000000000000000000000000001010"; -- 10
			op <= NOP;
			wait for clk_period;
			op <= ADDS;
			wait for clk_period;
			op <= ADDI;
			wait for clk_period;
			op <= SUBS;
			wait for clk_period;
			op <= SUBI;
			wait for clk_period;
			op <= ADDU;
			wait for clk_period;
			op <= ADDUI;
			wait for clk_period;
			op <= SUBU;
			wait for clk_period;
			op <= SUBUI;
			wait for clk_period;
			op <= ANDS;
			wait for clk_period;
			op <= ANDI;
			wait for clk_period;
			op <= ORS;
			wait for clk_period;
			op <= ORI;
			wait for clk_period;
			op <= XORS;
			wait for clk_period;
			op <= XORI;
			wait for clk_period;			
			op <= SEQI;
			wait for clk_period;
			op <= SNE;
			wait for clk_period;
			op <= SNEI;
			wait for clk_period;
			op <= SGEU;
			wait for clk_period;
			op <= SGEUI;
			wait for clk_period;
			op <= SLEU;
			wait for clk_period;
			op <= SLEUI;
			wait for clk_period;
			op <= SGTU;
			wait for clk_period;
			op <= SGTUI;
			wait for clk_period;			
			op <= SLTU;
			wait for clk_period;
			op <= SLTUI;
			wait for clk_period;
			op <= SGE;
			wait for clk_period;
			op <= SGEI;
			wait for clk_period;
			op <= SLE;
			wait for clk_period;
			op <= SLEI;
			wait for clk_period;
			op <= SGT;
			wait for clk_period;
			op <= SGTI;
			wait for clk_period;
			op <= SLTI;
			wait for clk_period;
			op <= SRLI;
			wait for clk_period;			
			op <= SLLS;
			wait for clk_period;
			op <= SLLI;
			wait for clk_period;
			op <= SRAS;
			wait for clk_period;
			op <= SRAI;
			wait for clk_period;
			in_A <= "00000000000000000000000000001010"; -- 10
			in_B <= "00000000000000000000000000110010"; -- 50
			op <= NOP;
			wait for clk_period;
			op <= ADDS;
			wait for clk_period;
			op <= ADDI;
			wait for clk_period;
			op <= SUBS;
			wait for clk_period;
			op <= SUBI;
			wait for clk_period;
			op <= ADDU;
			wait for clk_period;
			op <= ADDUI;
			wait for clk_period;
			op <= SUBU;
			wait for clk_period;
			op <= SUBUI;
			wait for clk_period;
			op <= ANDS;
			wait for clk_period;
			op <= ANDI;
			wait for clk_period;
			op <= ORS;
			wait for clk_period;
			op <= ORI;
			wait for clk_period;
			op <= XORS;
			wait for clk_period;
			op <= XORI;
			wait for clk_period;			
			op <= SEQI;
			wait for clk_period;
			op <= SNE;
			wait for clk_period;
			op <= SNEI;
			wait for clk_period;
			op <= SGEU;
			wait for clk_period;
			op <= SGEUI;
			wait for clk_period;
			op <= SLEU;
			wait for clk_period;
			op <= SLEUI;
			wait for clk_period;
			op <= SGTU;
			wait for clk_period;
			op <= SGTUI;
			wait for clk_period;			
			op <= SLTU;
			wait for clk_period;
			op <= SLTUI;
			wait for clk_period;
			op <= SGE;
			wait for clk_period;
			op <= SGEI;
			wait for clk_period;
			op <= SLE;
			wait for clk_period;
			op <= SLEI;
			wait for clk_period;
			op <= SGT;
			wait for clk_period;
			op <= SGTI;
			wait for clk_period;
			op <= SLTI;
			wait for clk_period;
			op <= SRLI;
			wait for clk_period;			
			op <= SLLS;
			wait for clk_period;
			op <= SLLI;
			wait for clk_period;
			op <= SRAS;
			wait for clk_period;
			op <= SRAI;
			wait for clk_period;
			in_A <= "00000000000000000000000000110010"; -- 50
			in_B <= "00000000000000000000000000001010"; -- 10
			op <= NOP;
			wait for clk_period;
			op <= ADDS;
			wait for clk_period;
			op <= ADDI;
			wait for clk_period;
			op <= SUBS;
			wait for clk_period;
			op <= SUBI;
			wait for clk_period;
			op <= ADDU;
			wait for clk_period;
			op <= ADDUI;
			wait for clk_period;
			op <= SUBU;
			wait for clk_period;
			op <= SUBUI;
			wait for clk_period;
			op <= ANDS;
			wait for clk_period;
			op <= ANDI;
			wait for clk_period;
			op <= ORS;
			wait for clk_period;
			op <= ORI;
			wait for clk_period;
			op <= XORS;
			wait for clk_period;
			op <= XORI;
			wait for clk_period;			
			op <= SEQI;
			wait for clk_period;
			op <= SNE;
			wait for clk_period;
			op <= SNEI;
			wait for clk_period;
			op <= SGEU;
			wait for clk_period;
			op <= SGEUI;
			wait for clk_period;
			op <= SLEU;
			wait for clk_period;
			op <= SLEUI;
			wait for clk_period;
			op <= SGTU;
			wait for clk_period;
			op <= SGTUI;
			wait for clk_period;			
			op <= SLTU;
			wait for clk_period;
			op <= SLTUI;
			wait for clk_period;
			op <= SGE;
			wait for clk_period;
			op <= SGEI;
			wait for clk_period;
			op <= SLE;
			wait for clk_period;
			op <= SLEI;
			wait for clk_period;
			op <= SGT;
			wait for clk_period;
			op <= SGTI;
			wait for clk_period;
			op <= SLTI;
			wait for clk_period;
			op <= SRLI;
			wait for clk_period;			
			op <= SLLS;
			wait for clk_period;
			op <= SLLI;
			wait for clk_period;
			op <= SRAS;
			wait for clk_period;
			op <= SRAI;
			wait for clk_period;
			in_A <= "11111111111111111111111111001110"; -- -50
			in_B <= "00000000000000000000000000001010"; -- 10
			op <= NOP;
			wait for clk_period;
			op <= ADDS;
			wait for clk_period;
			op <= ADDI;
			wait for clk_period;
			op <= SUBS;
			wait for clk_period;
			op <= SUBI;
			wait for clk_period;
			op <= ADDU;
			wait for clk_period;
			op <= ADDUI;
			wait for clk_period;
			op <= SUBU;
			wait for clk_period;
			op <= SUBUI;
			wait for clk_period;
			op <= ANDS;
			wait for clk_period;
			op <= ANDI;
			wait for clk_period;
			op <= ORS;
			wait for clk_period;
			op <= ORI;
			wait for clk_period;
			op <= XORS;
			wait for clk_period;
			op <= XORI;
			wait for clk_period;			
			op <= SEQI;
			wait for clk_period;
			op <= SNE;
			wait for clk_period;
			op <= SNEI;
			wait for clk_period;
			op <= SGEU;
			wait for clk_period;
			op <= SGEUI;
			wait for clk_period;
			op <= SLEU;
			wait for clk_period;
			op <= SLEUI;
			wait for clk_period;
			op <= SGTU;
			wait for clk_period;
			op <= SGTUI;
			wait for clk_period;			
			op <= SLTU;
			wait for clk_period;
			op <= SLTUI;
			wait for clk_period;
			op <= SGE;
			wait for clk_period;
			op <= SGEI;
			wait for clk_period;
			op <= SLE;
			wait for clk_period;
			op <= SLEI;
			wait for clk_period;
			op <= SGT;
			wait for clk_period;
			op <= SGTI;
			wait for clk_period;
			op <= SLTI;
			wait for clk_period;
			op <= SRLI;
			wait for clk_period;			
			op <= SLLS;
			wait for clk_period;
			op <= SLLI;
			wait for clk_period;
			op <= SRAS;
			wait for clk_period;
			op <= SRAI;
			wait for clk_period;			
			in_A <= "00000000000000000000000000001010"; -- 10
			in_B <= "11111111111111111111111111001110"; -- -50
			op <= NOP;
			wait for clk_period;
			op <= ADDS;
			wait for clk_period;
			op <= ADDI;
			wait for clk_period;
			op <= SUBS;
			wait for clk_period;
			op <= SUBI;
			wait for clk_period;
			op <= ADDU;
			wait for clk_period;
			op <= ADDUI;
			wait for clk_period;
			op <= SUBU;
			wait for clk_period;
			op <= SUBUI;
			wait for clk_period;
			op <= ANDS;
			wait for clk_period;
			op <= ANDI;
			wait for clk_period;
			op <= ORS;
			wait for clk_period;
			op <= ORI;
			wait for clk_period;
			op <= XORS;
			wait for clk_period;
			op <= XORI;
			wait for clk_period;			
			op <= SEQI;
			wait for clk_period;
			op <= SNE;
			wait for clk_period;
			op <= SNEI;
			wait for clk_period;
			op <= SGEU;
			wait for clk_period;
			op <= SGEUI;
			wait for clk_period;
			op <= SLEU;
			wait for clk_period;
			op <= SLEUI;
			wait for clk_period;
			op <= SGTU;
			wait for clk_period;
			op <= SGTUI;
			wait for clk_period;			
			op <= SLTU;
			wait for clk_period;
			op <= SLTUI;
			wait for clk_period;
			op <= SGE;
			wait for clk_period;
			op <= SGEI;
			wait for clk_period;
			op <= SLE;
			wait for clk_period;
			op <= SLEI;
			wait for clk_period;
			op <= SGT;
			wait for clk_period;
			op <= SGTI;
			wait for clk_period;
			op <= SLTI;
			wait for clk_period;
			op <= SRLI;
			wait for clk_period;			
			op <= SLLS;
			wait for clk_period;
			op <= SLLI;
			wait for clk_period;
			op <= SRAS;
			wait for clk_period;
			op <= SRAI;
			wait for clk_period;
			in_A <= "11111111111111111111111111110110"; -- -10
			in_B <= "11111111111111111111111111001110"; -- -50
			op <= NOP;
			wait for clk_period;
			op <= ADDS;
			wait for clk_period;
			op <= ADDI;
			wait for clk_period;
			op <= SUBS;
			wait for clk_period;
			op <= SUBI;
			wait for clk_period;
			op <= ADDU;
			wait for clk_period;
			op <= ADDUI;
			wait for clk_period;
			op <= SUBU;
			wait for clk_period;
			op <= SUBUI;
			wait for clk_period;
			op <= ANDS;
			wait for clk_period;
			op <= ANDI;
			wait for clk_period;
			op <= ORS;
			wait for clk_period;
			op <= ORI;
			wait for clk_period;
			op <= XORS;
			wait for clk_period;
			op <= XORI;
			wait for clk_period;			
			op <= SEQI;
			wait for clk_period;
			op <= SNE;
			wait for clk_period;
			op <= SNEI;
			wait for clk_period;
			op <= SGEU;
			wait for clk_period;
			op <= SGEUI;
			wait for clk_period;
			op <= SLEU;
			wait for clk_period;
			op <= SLEUI;
			wait for clk_period;
			op <= SGTU;
			wait for clk_period;
			op <= SGTUI;
			wait for clk_period;			
			op <= SLTU;
			wait for clk_period;
			op <= SLTUI;
			wait for clk_period;
			op <= SGE;
			wait for clk_period;
			op <= SGEI;
			wait for clk_period;
			op <= SLE;
			wait for clk_period;
			op <= SLEI;
			wait for clk_period;
			op <= SGT;
			wait for clk_period;
			op <= SGTI;
			wait for clk_period;
			op <= SLTI;
			wait for clk_period;
			op <= SRLI;
			wait for clk_period;			
			op <= SLLS;
			wait for clk_period;
			op <= SLLI;
			wait for clk_period;
			op <= SRAS;
			wait for clk_period;
			op <= SRAI;
			wait for clk_period;
			in_A <= "11111111111111111111111111001110"; -- -50
			in_B <= "11111111111111111111111111110110"; -- -10
			op <= NOP;
			wait for clk_period;
			op <= ADDS;
			wait for clk_period;
			op <= ADDI;
			wait for clk_period;
			op <= SUBS;
			wait for clk_period;
			op <= SUBI;
			wait for clk_period;
			op <= ADDU;
			wait for clk_period;
			op <= ADDUI;
			wait for clk_period;
			op <= SUBU;
			wait for clk_period;
			op <= SUBUI;
			wait for clk_period;
			op <= ANDS;
			wait for clk_period;
			op <= ANDI;
			wait for clk_period;
			op <= ORS;
			wait for clk_period;
			op <= ORI;
			wait for clk_period;
			op <= XORS;
			wait for clk_period;
			op <= XORI;
			wait for clk_period;			
			op <= SEQI;
			wait for clk_period;
			op <= SNE;
			wait for clk_period;
			op <= SNEI;
			wait for clk_period;
			op <= SGEU;
			wait for clk_period;
			op <= SGEUI;
			wait for clk_period;
			op <= SLEU;
			wait for clk_period;
			op <= SLEUI;
			wait for clk_period;
			op <= SGTU;
			wait for clk_period;
			op <= SGTUI;
			wait for clk_period;			
			op <= SLTU;
			wait for clk_period;
			op <= SLTUI;
			wait for clk_period;
			op <= SGE;
			wait for clk_period;
			op <= SGEI;
			wait for clk_period;
			op <= SLE;
			wait for clk_period;
			op <= SLEI;
			wait for clk_period;
			op <= SGT;
			wait for clk_period;
			op <= SGTI;
			wait for clk_period;
			op <= SLTI;
			wait for clk_period;
			op <= SRLI;
			wait for clk_period;			
			op <= SLLS;
			wait for clk_period;
			op <= SLLI;
			wait for clk_period;
			op <= SRAS;
			wait for clk_period;
			op <= SRAI;
			wait for clk_period;			
			in_A <= "11111111111111111111111111110110"; -- -10
			in_B <= "11111111111111111111111111110110"; -- -10
			op <= NOP;
			wait for clk_period;
			op <= ADDS;
			wait for clk_period;
			op <= ADDI;
			wait for clk_period;
			op <= SUBS;
			wait for clk_period;
			op <= SUBI;
			wait for clk_period;
			op <= ADDU;
			wait for clk_period;
			op <= ADDUI;
			wait for clk_period;
			op <= SUBU;
			wait for clk_period;
			op <= SUBUI;
			wait for clk_period;
			op <= ANDS;
			wait for clk_period;
			op <= ANDI;
			wait for clk_period;
			op <= ORS;
			wait for clk_period;
			op <= ORI;
			wait for clk_period;
			op <= XORS;
			wait for clk_period;
			op <= XORI;
			wait for clk_period;			
			op <= SEQI;
			wait for clk_period;
			op <= SNE;
			wait for clk_period;
			op <= SNEI;
			wait for clk_period;
			op <= SGEU;
			wait for clk_period;
			op <= SGEUI;
			wait for clk_period;
			op <= SLEU;
			wait for clk_period;
			op <= SLEUI;
			wait for clk_period;
			op <= SGTU;
			wait for clk_period;
			op <= SGTUI;
			wait for clk_period;			
			op <= SLTU;
			wait for clk_period;
			op <= SLTUI;
			wait for clk_period;
			op <= SGE;
			wait for clk_period;
			op <= SGEI;
			wait for clk_period;
			op <= SLE;
			wait for clk_period;
			op <= SLEI;
			wait for clk_period;
			op <= SGT;
			wait for clk_period;
			op <= SGTI;
			wait for clk_period;
			op <= SLTI;
			wait for clk_period;
			op <= SRLI;
			wait for clk_period;			
			op <= SLLS;
			wait for clk_period;
			op <= SLLI;
			wait for clk_period;
			op <= SRAS;
			wait for clk_period;
			op <= SRAI;
			wait for clk_period;
			in_A <= "00000000000000000000000000000000"; -- 0
			in_B <= "11111111111111111111111111110110"; -- -10
			op <= NOP;
			wait for clk_period;
			op <= ADDS;
			wait for clk_period;
			op <= ADDI;
			wait for clk_period;
			op <= SUBS;
			wait for clk_period;
			op <= SUBI;
			wait for clk_period;
			op <= ADDU;
			wait for clk_period;
			op <= ADDUI;
			wait for clk_period;
			op <= SUBU;
			wait for clk_period;
			op <= SUBUI;
			wait for clk_period;
			op <= ANDS;
			wait for clk_period;
			op <= ANDI;
			wait for clk_period;
			op <= ORS;
			wait for clk_period;
			op <= ORI;
			wait for clk_period;
			op <= XORS;
			wait for clk_period;
			op <= XORI;
			wait for clk_period;			
			op <= SEQI;
			wait for clk_period;
			op <= SNE;
			wait for clk_period;
			op <= SNEI;
			wait for clk_period;
			op <= SGEU;
			wait for clk_period;
			op <= SGEUI;
			wait for clk_period;
			op <= SLEU;
			wait for clk_period;
			op <= SLEUI;
			wait for clk_period;
			op <= SGTU;
			wait for clk_period;
			op <= SGTUI;
			wait for clk_period;			
			op <= SLTU;
			wait for clk_period;
			op <= SLTUI;
			wait for clk_period;
			op <= SGE;
			wait for clk_period;
			op <= SGEI;
			wait for clk_period;
			op <= SLE;
			wait for clk_period;
			op <= SLEI;
			wait for clk_period;
			op <= SGT;
			wait for clk_period;
			op <= SGTI;
			wait for clk_period;
			op <= SLTI;
			wait for clk_period;
			op <= SRLI;
			wait for clk_period;			
			op <= SLLS;
			wait for clk_period;
			op <= SLLI;
			wait for clk_period;
			op <= SRAS;
			wait for clk_period;
			op <= SRAI;
			wait for clk_period;
			in_A <= "11111111111111111111111111110110"; -- -10
			in_B <= "00000000000000000000000000000000"; -- 0			
			op <= NOP;
			wait for clk_period;
			op <= ADDS;
			wait for clk_period;
			op <= ADDI;
			wait for clk_period;
			op <= SUBS;
			wait for clk_period;
			op <= SUBI;
			wait for clk_period;
			op <= ADDU;
			wait for clk_period;
			op <= ADDUI;
			wait for clk_period;
			op <= SUBU;
			wait for clk_period;
			op <= SUBUI;
			wait for clk_period;
			op <= ANDS;
			wait for clk_period;
			op <= ANDI;
			wait for clk_period;
			op <= ORS;
			wait for clk_period;
			op <= ORI;
			wait for clk_period;
			op <= XORS;
			wait for clk_period;
			op <= XORI;
			wait for clk_period;			
			op <= SEQI;
			wait for clk_period;
			op <= SNE;
			wait for clk_period;
			op <= SNEI;
			wait for clk_period;
			op <= SGEU;
			wait for clk_period;
			op <= SGEUI;
			wait for clk_period;
			op <= SLEU;
			wait for clk_period;
			op <= SLEUI;
			wait for clk_period;
			op <= SGTU;
			wait for clk_period;
			op <= SGTUI;
			wait for clk_period;			
			op <= SLTU;
			wait for clk_period;
			op <= SLTUI;
			wait for clk_period;
			op <= SGE;
			wait for clk_period;
			op <= SGEI;
			wait for clk_period;
			op <= SLE;
			wait for clk_period;
			op <= SLEI;
			wait for clk_period;
			op <= SGT;
			wait for clk_period;
			op <= SGTI;
			wait for clk_period;
			op <= SLTI;
			wait for clk_period;
			op <= SRLI;
			wait for clk_period;			
			op <= SLLS;
			wait for clk_period;
			op <= SLLI;
			wait for clk_period;
			op <= SRAS;
			wait for clk_period;
			op <= SRAI;
			wait for clk_period;	
			in_A <= "00000000000000000000000000000000"; -- 0
			in_B <= "00000000000000000000000000000000"; -- 0			
			op <= NOP;
			wait for clk_period;
			op <= ADDS;
			wait for clk_period;
			op <= ADDI;
			wait for clk_period;
			op <= SUBS;
			wait for clk_period;
			op <= SUBI;
			wait for clk_period;
			op <= ADDU;
			wait for clk_period;
			op <= ADDUI;
			wait for clk_period;
			op <= SUBU;
			wait for clk_period;
			op <= SUBUI;
			wait for clk_period;
			op <= ANDS;
			wait for clk_period;
			op <= ANDI;
			wait for clk_period;
			op <= ORS;
			wait for clk_period;
			op <= ORI;
			wait for clk_period;
			op <= XORS;
			wait for clk_period;
			op <= XORI;
			wait for clk_period;			
			op <= SEQI;
			wait for clk_period;
			op <= SNE;
			wait for clk_period;
			op <= SNEI;
			wait for clk_period;
			op <= SGEU;
			wait for clk_period;
			op <= SGEUI;
			wait for clk_period;
			op <= SLEU;
			wait for clk_period;
			op <= SLEUI;
			wait for clk_period;
			op <= SGTU;
			wait for clk_period;
			op <= SGTUI;
			wait for clk_period;			
			op <= SLTU;
			wait for clk_period;
			op <= SLTUI;
			wait for clk_period;
			op <= SGE;
			wait for clk_period;
			op <= SGEI;
			wait for clk_period;
			op <= SLE;
			wait for clk_period;
			op <= SLEI;
			wait for clk_period;
			op <= SGT;
			wait for clk_period;
			op <= SGTI;
			wait for clk_period;
			op <= SLTI;
			wait for clk_period;
			op <= SRLI;
			wait for clk_period;			
			op <= SLLS;
			wait for clk_period;
			op <= SLLI;
			wait for clk_period;
			op <= SRAS;
			wait for clk_period;
			op <= SRAI;
			wait for clk_period;
	end process;
end architecture test;	